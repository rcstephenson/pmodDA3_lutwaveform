-- Ryan Stephenson jan 20 2020
-- welcome to my little slice of memory :)
-- 01/24 updated to 41 datapoints for 25MHz clock  
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is 
    generic( N : integer := 7; --array length = 2**N
             M : integer := 16); --data width
    port(
         clk : in std_logic;
        ADDR : in std_logic_vector(N-1 downto 0);
          en : in std_logic; --active low
        Dout : out std_logic_vector(M-1 downto 0)
    );
end ROM;

architecture behv of ROM is 
    type ROM is array(0 to 82-1) of std_logic_vector(M-1 downto 0); 
    signal mem : ROM := ("0000000000000000", "0000000110010100", "0000001100101001", "0000010010111101", "0000011001010010", "0000011111100110", "0000100101111011", "0000101100001111", "0000110010100100", "0000111000111000", "0000111111001101", "0001000101100001", "0001001011110110", "0001010010001010", "0001011000011111", "0001011110110011", "0001100101001000", "0001101011011101", "0001110001110001", "0001111000000110", "0001111110011010", "0010000100101111", "0010001011000011", "0010010001011000", "0010010111101100", "0010011110000001", "0010100100010101", "0010101010101010", "0010110000111110", "0010110111010011", "0010111101100111", "0011000011111100", "0011001010010000", "0011010000100101", "0011010110111010", "0011011101001110", "0011100011100011", "0011101001110111", "0011110000001100", "0011110110100000", "0011111100110101", "0100000011001001", "0100001001011110", "0100001111110010", "0100010110000111", "0100011100011011", "0100100010110000", "0100101001000100", "0100101111011001", "0100110101101110", "0100111100000010", "0101000010010111", "0101001000101011", "0101001111000000", "0101010101010100", "0101011011101001", "0101100001111101", "0101101000010010", "0101101110100110", "0101110100111011", "0101111011001111", "0110000001100100", "0110000111111000", "0110001110001101", "0110010100100001", "0110011010110110", "0110100001001011", "0110100111011111", "0110101101110100", "0110110100001000", "0110111010011101", "0111000000110001", "0111000111000110", "0111001101011010", "0111010011101111", "0111011010000011", "0111100000011000", "0111100110101100", "0111101101000001", "0111110011010101", "0111111001101010", "0111111111111111");
        begin 
    process(clk,en,ADDR)
    begin 
        if (clk'event and clk='1') then 
            if (en='0') then --D_out logic
                Dout <= mem(to_integer(unsigned(ADDR)));
            else
                Dout <= (others => '0');
            end if;
        end if;
    end process;
end behv;